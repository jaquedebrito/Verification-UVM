//------------------------------------------------------------------------------
// File: sqrt_test_pkg.sv
// Author: Jaqueline F. de Brito
// Date: 2025-03-28 17:10:24
//------------------------------------------------------------------------------

`include "uvm_macros.svh"
`include "bvm_macros.svh"

package sqrt_test_pkg;

    import uvm_pkg::*;
    import bvm_pkg::*;

    `include "sqrt_transaction.svh"
    `include "sqrt_sequence.svh"
    typedef uvm_sequencer #(sqrt_transaction) sqrt_sequencer;
    `include "sqrt_driver.svh"
    `include "sqrt_monitor.svh"
    `include "sqrt_agent.svh"
    `include "sqrt_coverage_in.svh"
    `include "sqrt_coverage_out.svh"
    `include "sqrt_refmod.svh"
    `include "sqrt_env.svh"
    `include "sqrt_test.svh"

endpackage